// bypass multiplexer
`define HZ_BYPASS_NONE 2'b00
`define HZ_BYPASS_W2E  2'b01
`define HZ_BYPASS_M2E  2'b10
