`define LDST_B      3'd0    // signed  byte
`define LDST_H      3'd1    // signed  half-world
`define LDST_W      3'd2    // word
`define LDST_BU     3'd4    // unsigned byte (only for read)
`define LDST_HU     3'd5    // unsigned half-world (only for read)